LIBRARY ieee;
USE ieee.STD_LOGIC_1164.all;

ENTITY two_one_multi IS 
  PORT(
       SW:IN STD_LOGIC_VECTOR(17 DOWNTO 0 );
       LEDR: OUT STD_LOGIC_VECTOR(17 DOWNTO 0);
       LEDG: OUT STD_LOGIC_VECTOR(17 DOWNTO 0);
       m:BUFFER STD_LOGIC_VECTOR(7 DOWNTO 0));
END two_one_multi;

ARCHITECTURE Behavior OF two_one_multi IS

BEGIN
  

  WITH SW(17 DOWNTO 1) SELECT
  m<= SW(7 DOWNTO 0) WHEN '0',
      SW(15 DOWNTO 8) WHEN '1',
      "00000000" WHEN OTHERS;


  LEDR <= SW;
  LEDG(7 DOWNTO 0) <= m;
END Behavior;






