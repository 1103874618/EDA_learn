LIBRARY ieee;
USE ieee.STD_LOGIC_1164.all;

ENTITY seven_segment_decoder IS 
PORT(
       HEX0: OUT STD_LOGIC_VECTOR(0 TO 6);--0为灯亮
       SW:IN STD_LOGIC_VECTOR(17 DOWNTO 0 );
       LEDR: OUT STD_LOGIC_VECTOR(17 DOWNTO 0);
       LEDG: OUT STD_LOGIC_VECTOR(17 DOWNTO 0));
END seven_segment_decoder;

ARCHITECTURE Behavior OF seven_segment_decoder IS
BEGIN

HEX0<="1001000" WHEN SW(2 DOWNTO 1)="00" ELSE
      "0110000" WHEN SW(2 DOWNTO 1)="01" ELSE
      "1110001" WHEN SW(2 DOWNTO 1)="10" ELSE
      "0000001" WHEN SW(2 DOWNTO 1)="11" ELSE
      "1111111";

END Behavior;



